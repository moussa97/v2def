
VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS DATABASE MICRONS 1000 ;
END UNITS

USEMINSPACING OBS ON ;
USEMINSPACING PIN OFF ;
CLEARANCEMEASURE EUCLIDEAN ;


MANUFACTURINGGRID 0.1 ;

LAYER nwell
  TYPE	MASTERSLICE ;
END nwell

LAYER nactive
  TYPE	MASTERSLICE ;
END nactive

LAYER pactive
  TYPE	MASTERSLICE ;
END pactive

LAYER poly
  TYPE	MASTERSLICE ;
END poly

LAYER cc
  TYPE	CUT ;
  SPACING	0.9 ;
END cc

LAYER metal1
  TYPE		ROUTING ;
  DIRECTION	HORIZONTAL ;
  PITCH		2  ;
  WIDTH		0.6 ;
  SPACING	0.6 ;
  OFFSET	1 ;
  RESISTANCE	RPERSQ 0.07 ;
  CAPACITANCE	CPERSQDIST 3e-05 ;
END metal1

LAYER via1
  TYPE	CUT ;
  SPACING	0.6 ;
END via1



VIA M2_M1 DEFAULT
  LAYER metal1 ;
    RECT -0.400 -0.400 0.400 0.400 ;
  LAYER via1 ;
    RECT -0.200 -0.200 0.200 0.200 ;
  LAYER metal2 ;
    RECT -0.400 -0.400 0.400 0.400 ;
END M2_M1

VIA M3_M2 DEFAULT
  LAYER metal2 ;
    RECT -0.400 -0.400 0.400 0.400 ;
  LAYER via2 ;
    RECT -0.200 -0.200 0.200 0.200 ;
  LAYER metal3 ;
    RECT -0.400 -0.400 0.400 0.400 ;
END M3_M2