
VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS DATABASE MICRONS 1000 ;
END UNITS

USEMINSPACING OBS ON ;
USEMINSPACING PIN OFF ;
CLEARANCEMEASURE EUCLIDEAN ;


MANUFACTURINGGRID 0.1 ;

LAYER nwell
  TYPE	MASTERSLICE ;
END nwell

LAYER nactive
  TYPE	MASTERSLICE ;
END nactive

LAYER pactive
  TYPE	MASTERSLICE ;
END pactive

LAYER poly
  TYPE	MASTERSLICE ;
END poly

LAYER cc
  TYPE	CUT ;
  SPACING	0.9 ;
END cc

LAYER metal1
  TYPE		ROUTING ;
  DIRECTION	HORIZONTAL ;
  PITCH		2  ;
  WIDTH		0.6 ;
  SPACING	0.6 ;
  OFFSET	1 ;
  RESISTANCE	RPERSQ 0.07 ;
  CAPACITANCE	CPERSQDIST 3e-05 ;
END metal1

LAYER via1

  TYPE	CUT ;
  SPACING	0.6 ;
END via1

LAYER metal2
  TYPE		ROUTING ;
  DIRECTION	VERTICAL ;
  PITCH		1.6  ;
  WIDTH		0.6 ;
  SPACING	0.6 ;
  OFFSET	0.8 ;
  RESISTANCE	RPERSQ 0.07 ;
  CAPACITANCE	CPERSQDIST 1.7e-05 ;
END metal2

LAYER via2
  TYPE	CUT ;
  SPACING	0.6 ;
END via2

LAYER metal3
  TYPE		ROUTING ;
  DIRECTION	HORIZONTAL ;
  PITCH		2  ;
  WIDTH		0.6 ;
  SPACING	0.6 ;
  OFFSET	1 ;
  RESISTANCE	RPERSQ 0.07 ;
  CAPACITANCE	CPERSQDIST 7e-06 ;
END metal3

LAYER via3
  TYPE	CUT ;
  SPACING	0.8 ;
END via3

LAYER metal4
  TYPE		ROUTING ;
  DIRECTION	VERTICAL ;
  PITCH		3.2  ;
  WIDTH		1.2 ;
  SPACING	1.2 ;
  OFFSET	1.6 ;
  RESISTANCE	RPERSQ 0.04 ;
  CAPACITANCE	CPERSQDIST 4e-06 ;
END metal4

VIA M2_M1 DEFAULT
  LAYER metal1 ;
    RECT -0.400 -0.400 0.400 0.400 ;
  LAYER via1 ;
    RECT -0.200 -0.200 0.200 0.200 ;
  LAYER metal2 ;
    RECT -0.400 -0.400 0.400 0.400 ;
END M2_M1

VIA M3_M2 DEFAULT
  LAYER metal2 ;
    RECT -0.400 -0.400 0.400 0.400 ;
  LAYER via2 ;
    RECT -0.200 -0.200 0.200 0.200 ;
  LAYER metal3 ;
    RECT -0.400 -0.400 0.400 0.400 ;
END M3_M2

VIA M4_M3 DEFAULT
  LAYER metal3 ;
    RECT -0.400 -0.400 0.400 0.400 ;
  LAYER via3 ;
    RECT -0.200 -0.200 0.200 0.200 ;
  LAYER metal4 ;
    RECT -0.600 -0.600 0.600 0.600 ;
END M4_M3


SITE  corner
    CLASS	PAD ;
    SYMMETRY	R90 Y ;
    SIZE	300.000 BY 300.000 ;
END  corner

SITE  IO
    CLASS	PAD ;
    SYMMETRY	Y ;
    SIZE	90.000 BY 300.000 ;
END  IO

SITE  core
    CLASS	CORE ;
    SYMMETRY	Y ;
    SIZE	1.600 BY 20.000 ;
END  core

MACRO FILL
  CLASS  CORE ;
  FOREIGN FILL 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.600 BY 20.000 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.400 -0.600 2.000 0.600 ;
    END
  END gnd
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.400 19.400 2.000 20.600 ;
    END
  END vdd
END FILL

MACRO AND2X1
  CLASS  CORE ;
  FOREIGN AND2X1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.400 BY 20.000 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
	
    PORT
      LAYER metal1 ;
        RECT 0.400 6.600 1.200 8.200 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        RECT 2.600 9.800 3.400 11.400 ;
        RECT 2.000 10.600 3.400 11.400 ;
    END
  END B
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 3.000 -0.600 3.800 5.200 ;
        RECT -0.400 -0.600 6.800 0.600 ;
    END
  END gnd
  PIN Y
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        RECT 5.200 12.600 6.000 13.400 ;
        RECT 5.200 14.800 6.000 18.800 ;
        RECT 5.400 3.200 6.000 18.800 ;
        RECT 4.600 1.200 5.400 3.800 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.400 14.800 1.200 20.600 ;
        RECT -0.400 19.400 6.800 20.600 ;
        RECT 3.600 14.800 4.400 20.600 ;
    END
  END vdd
  OBS 
      LAYER metal1 ;
        RECT 0.400 1.200 1.200 5.200 ;
        RECT 0.600 5.200 2.400 5.800 ;
        RECT 1.800 5.200 2.400 6.600 ;
        RECT 4.000 5.800 4.800 6.600 ;
        RECT 1.800 6.000 4.800 6.600 ;
        RECT 4.000 5.800 4.600 14.200 ;
        RECT 2.200 13.600 4.600 14.200 ;
        RECT 2.200 13.600 2.800 18.800 ;
        RECT 2.000 14.800 2.800 18.800 ;
  END 
END AND2X1

MACRO AND2X2
  CLASS  CORE ;
  FOREIGN AND2X2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.400 BY 20.000 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        RECT 0.400 6.600 1.200 8.200 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        RECT 2.200 7.200 2.800 9.400 ;
        RECT 2.400 7.000 3.200 7.800 ;
        RECT 2.000 8.600 2.800 9.400 ;
    END
  END B
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 3.000 -0.600 3.800 5.000 ;
        RECT -0.400 -0.600 6.800 0.600 ;
    END
  END gnd
  PIN Y
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        RECT 5.200 8.600 6.000 9.400 ;
        RECT 5.200 10.800 6.000 18.800 ;
        RECT 5.400 4.200 6.000 18.800 ;
        RECT 4.600 1.200 5.400 5.200 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.400 14.800 1.200 20.600 ;
        RECT -0.400 19.400 6.800 20.600 ;
        RECT 3.600 11.200 4.400 20.600 ;
    END
  END vdd
  OBS 
      LAYER metal1 ;
        RECT 0.400 1.200 1.200 5.200 ;
        RECT 0.600 1.200 1.200 6.000 ;
        RECT 0.600 5.400 2.400 6.000 ;
        RECT 1.800 5.800 4.800 6.400 ;
        RECT 4.000 5.800 4.800 6.600 ;
        RECT 4.000 5.800 4.600 10.600 ;
        RECT 2.200 10.000 4.600 10.600 ;
        RECT 2.200 10.000 2.800 18.800 ;
        RECT 2.000 14.800 2.800 18.800 ;
  END 
END AND2X2

MACRO AOI21X1
  CLASS  CORE ;
  FOREIGN AOI21X1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.400 BY 20.000 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        RECT 0.400 8.600 1.200 9.400 ;
        RECT 1.200 8.800 2.000 9.800 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        RECT 2.000 6.600 2.800 8.200 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        RECT 5.000 3.800 5.800 4.600 ;
        RECT 5.200 4.600 6.000 5.400 ;
    END
  END C
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 1.000 -0.600 1.800 5.200 ;
        RECT -0.400 -0.600 6.800 0.600 ;
        RECT 5.200 -0.600 6.000 3.200 ;
    END
  END gnd
  PIN Y
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        RECT 3.600 1.200 4.200 9.400 ;
        RECT 5.200 10.800 6.000 18.800 ;
        RECT 3.600 8.800 6.000 9.400 ;
        RECT 5.200 8.600 6.000 9.400 ;
        RECT 5.200 8.600 5.800 18.800 ;
        RECT 3.600 1.200 4.400 5.200 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 2.000 12.000 2.800 20.600 ;
        RECT -0.400 19.400 6.800 20.600 ;
    END
  END vdd
  OBS 
      LAYER metal1 ;
        RECT 0.400 10.800 4.400 11.400 ;
        RECT 0.400 10.800 1.200 18.800 ;
        RECT 3.600 10.800 4.400 18.800 ;
  END 
END AOI21X1

MACRO AOI22X1
  CLASS  CORE ;
  FOREIGN AOI22X1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.000 BY 20.000 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        RECT 0.400 8.600 1.200 9.400 ;
        RECT 1.200 8.800 2.000 9.800 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        RECT 2.000 6.600 2.800 8.200 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        RECT 6.800 8.600 7.600 10.200 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        RECT 5.200 6.600 5.800 8.600 ;
        RECT 5.200 6.600 6.000 7.400 ;
        RECT 5.000 7.800 5.800 8.600 ;
    END
  END D
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.800 -0.600 1.600 5.200 ;
        RECT -0.400 -0.600 8.400 0.600 ;
        RECT 6.800 -0.600 7.600 5.200 ;
    END
  END gnd
  PIN Y
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        RECT 3.600 8.600 4.400 9.400 ;
        RECT 5.200 10.800 6.000 17.600 ;
        RECT 5.200 9.600 5.800 17.600 ;
        RECT 3.800 9.600 5.800 10.200 ;
        RECT 3.400 1.200 5.000 5.200 ;
        RECT 3.800 1.200 4.400 10.200 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 2.000 12.000 2.800 20.600 ;
        RECT -0.400 19.400 8.400 20.600 ;
    END
  END vdd
  OBS 
      LAYER metal1 ;
        RECT 0.400 10.800 4.400 11.400 ;
        RECT 3.600 10.800 4.400 18.800 ;
        RECT 0.400 10.800 1.200 18.800 ;
        RECT 6.800 10.800 7.600 18.800 ;
        RECT 3.600 18.200 7.600 18.800 ;
  END 
END AOI22X1

MACRO BUFX2
  CLASS  CORE ;
  FOREIGN BUFX2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.800 BY 20.000 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        RECT 0.400 7.800 1.200 9.400 ;
    END
  END A
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 2.000 -0.600 2.800 5.200 ;
        RECT -0.400 -0.600 5.200 0.600 ;
    END
  END gnd
  PIN Y
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        RECT 3.600 1.200 4.400 8.600 ;
        RECT 3.600 10.800 4.400 18.800 ;
        RECT 3.800 1.200 4.400 18.800 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 2.000 12.000 2.800 20.600 ;
        RECT -0.400 19.400 5.200 20.600 ;
    END
  END vdd
  OBS 
      LAYER metal1 ;
        RECT 0.400 1.200 1.200 6.400 ;
        RECT 0.400 5.800 2.600 6.400 ;
        RECT 2.000 9.400 3.200 10.200 ;
        RECT 2.000 5.800 2.600 11.400 ;
        RECT 0.400 10.800 2.600 11.400 ;
        RECT 0.400 10.800 1.200 18.800 ;
  END 
END BUFX2

MACRO BUFX4
  CLASS  CORE ;
  FOREIGN BUFX4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.400 BY 20.000 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        RECT 0.600 7.800 1.400 9.400 ;
        RECT 0.400 8.600 1.400 9.400 ;
    END
  END A
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 2.000 -0.600 2.800 5.200 ;
        RECT -0.400 -0.600 6.800 0.600 ;
        RECT 5.200 -0.600 6.000 5.200 ;
    END
  END gnd
  PIN Y
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        RECT 3.600 1.200 4.400 5.200 ;
        RECT 4.000 4.600 4.600 11.800 ;
        RECT 3.600 10.800 4.400 18.800 ;
        RECT 3.600 6.600 4.600 7.400 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 2.000 12.000 2.800 20.600 ;
        RECT -0.400 19.400 6.800 20.600 ;
        RECT 5.200 10.800 6.000 20.600 ;
    END
  END vdd
  OBS 
      LAYER metal1 ;
        RECT 0.400 1.200 1.200 6.400 ;
        RECT 0.400 5.800 3.000 6.400 ;
        RECT 2.400 8.000 3.400 8.800 ;
        RECT 2.400 5.800 3.000 11.400 ;
        RECT 0.400 10.800 3.000 11.400 ;
        RECT 0.400 10.800 1.200 18.800 ;
  END 
END BUFX4

MACRO DFFNEGX1
  CLASS  CORE ;
  FOREIGN DFFNEGX1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 19.200 BY 20.000 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        RECT 14.600 9.400 15.400 10.200 ;
        RECT 18.000 1.200 18.800 18.800 ;
        RECT 14.600 9.600 18.800 10.200 ;
        RECT 15.000 5.600 18.800 6.200 ;
        RECT 15.000 5.400 15.800 6.200 ;
    END
  END Q
  PIN CLK
    DIRECTION INPUT ;
    PORT
      LAYER metal2 ;
        RECT 5.200 6.800 6.000 13.400 ;
      LAYER via1 ;
        RECT 5.400 12.800 5.800 13.200 ;
        RECT 5.400 7.000 5.800 7.400 ;
      LAYER metal1 ;
        RECT 5.200 12.600 6.000 13.400 ;
        RECT 1.200 6.800 12.800 7.400 ;
        RECT 12.000 6.600 12.800 7.400 ;
        RECT 5.200 6.800 6.000 7.600 ;
        RECT 4.200 4.600 5.000 5.400 ;
        RECT 4.000 5.400 4.800 7.400 ;
        RECT 1.200 6.600 2.800 7.400 ;
        RECT 5.400 13.400 6.200 14.200 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        RECT 2.800 8.400 3.600 9.200 ;
        RECT 6.800 8.600 7.600 9.400 ;
        RECT 2.800 8.600 7.600 9.200 ;
    END
  END D
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 2.000 -0.600 2.800 5.200 ;
        RECT -0.400 -0.600 19.600 0.600 ;
        RECT 16.400 -0.600 17.200 5.000 ;
        RECT 10.800 -0.600 11.600 3.200 ;
        RECT 7.400 -0.600 8.400 3.200 ;
    END
  END gnd
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 2.000 11.000 2.800 20.600 ;
        RECT -0.400 19.400 19.600 20.600 ;
        RECT 16.400 10.800 17.200 20.600 ;
        RECT 10.800 14.800 11.600 20.600 ;
        RECT 7.600 14.800 8.400 20.600 ;
    END
  END vdd
  OBS 
      LAYER metal2 ;
        RECT 0.400 5.200 1.200 10.800 ;
        RECT 3.600 3.200 4.400 10.000 ;
        RECT 3.600 3.200 4.200 14.800 ;
        RECT 3.600 10.800 4.400 14.800 ;
        RECT 13.200 3.200 14.000 11.400 ;
        RECT 13.200 3.200 13.800 14.800 ;
        RECT 13.200 12.200 14.000 14.800 ;
      LAYER metal1 ;
        RECT 0.400 1.200 1.200 6.000 ;
        RECT 3.600 14.000 4.400 15.400 ;
        RECT 3.600 14.800 5.600 15.400 ;
        RECT 4.800 14.800 5.600 18.800 ;
        RECT 4.800 1.200 5.600 3.200 ;
        RECT 3.600 2.600 5.600 3.200 ;
        RECT 3.600 2.600 4.400 4.000 ;
        RECT 3.600 11.400 9.000 12.000 ;
        RECT 3.600 11.400 4.400 12.200 ;
        RECT 8.200 11.400 9.000 12.200 ;
        RECT 9.200 1.200 10.000 3.200 ;
        RECT 9.200 1.200 9.800 4.400 ;
        RECT 7.000 3.800 9.800 4.400 ;
        RECT 7.000 3.800 7.800 4.600 ;
        RECT 7.000 13.400 7.800 14.200 ;
        RECT 9.800 13.400 10.600 14.200 ;
        RECT 7.000 13.600 10.600 14.200 ;
        RECT 9.200 13.600 9.800 18.800 ;
        RECT 9.200 14.800 10.000 18.800 ;
        RECT 13.200 14.000 14.000 14.800 ;
        RECT 13.400 14.800 14.600 18.800 ;
        RECT 0.400 9.800 5.000 10.400 ;
        RECT 4.200 10.200 11.400 10.800 ;
        RECT 10.800 10.200 11.400 12.200 ;
        RECT 10.800 11.400 14.600 12.000 ;
        RECT 10.800 11.400 11.800 12.200 ;
        RECT 13.800 11.400 14.600 12.200 ;
        RECT 0.400 9.800 1.200 18.800 ;
        RECT 13.400 1.200 14.600 3.200 ;
        RECT 13.200 2.600 14.000 4.000 ;
        RECT 13.200 8.000 14.000 8.800 ;
        RECT 13.200 8.200 17.000 8.800 ;
        RECT 16.200 8.200 17.000 9.000 ;
      LAYER via1 ;
        RECT 0.600 10.200 1.000 10.600 ;
        RECT 0.600 5.400 1.000 5.800 ;
        RECT 3.800 14.200 4.200 14.600 ;
        RECT 3.800 11.600 4.200 12.000 ;
        RECT 3.800 3.400 4.200 3.800 ;
        RECT 13.400 14.200 13.800 14.600 ;
        RECT 13.400 8.200 13.800 8.600 ;
        RECT 13.400 3.400 13.800 3.800 ;
  END 
END DFFNEGX1

MACRO NOR3X1
  CLASS  CORE ;
  FOREIGN NOR3X1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.800 BY 20.000 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        RECT 2.000 4.600 3.800 5.400 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        RECT 3.600 6.600 5.200 7.400 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        RECT 5.200 8.600 6.800 9.400 ;
    END
  END C
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 2.000 -0.600 2.800 3.200 ;
        RECT -0.400 -0.600 13.200 0.600 ;
        RECT 5.200 -0.600 6.000 2.800 ;
    END
  END gnd
  PIN Y
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        RECT 3.600 1.200 4.400 3.200 ;
        RECT 10.000 12.000 10.800 17.600 ;
        RECT 10.000 10.600 10.800 11.400 ;
        RECT 10.000 10.600 10.600 17.600 ;
        RECT 7.400 10.600 10.800 11.200 ;
        RECT 7.400 3.200 8.000 11.200 ;
        RECT 6.800 1.200 7.600 4.000 ;
        RECT 4.000 3.400 8.000 4.000 ;
        RECT 4.000 2.600 4.600 4.000 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 2.000 12.800 2.800 20.600 ;
        RECT -0.400 19.400 13.200 20.600 ;
    END
  END vdd
  OBS 
      LAYER metal1 ;
        RECT 0.600 11.600 4.200 12.200 ;
        RECT 3.600 11.600 4.200 18.800 ;
        RECT 3.600 12.800 4.400 18.800 ;
        RECT 0.600 11.600 1.200 18.800 ;
        RECT 0.400 12.800 1.200 18.800 ;
        RECT 6.800 13.000 7.600 18.800 ;
        RECT 3.600 18.200 7.600 18.800 ;
        RECT 5.400 11.800 9.000 12.400 ;
        RECT 5.400 11.800 6.000 17.600 ;
        RECT 5.200 12.800 6.000 17.600 ;
        RECT 8.400 12.000 9.200 18.000 ;
        RECT 11.600 12.000 12.400 18.000 ;
        RECT 8.600 12.000 9.200 18.800 ;
        RECT 11.600 12.000 12.200 18.800 ;
        RECT 8.600 18.200 12.200 18.800 ;
  END 
END NOR3X1

MACRO DFFPOSX1
  CLASS  CORE ;
  FOREIGN DFFPOSX1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 19.200 BY 20.000 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        RECT 14.600 9.400 15.400 10.200 ;
        RECT 18.000 1.200 18.800 18.800 ;
        RECT 14.600 9.600 18.800 10.200 ;
        RECT 15.000 5.600 18.800 6.200 ;
        RECT 15.000 5.400 15.800 6.200 ;
    END
  END Q
  PIN CLK
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        RECT 1.200 6.600 2.800 7.400 ;
        RECT 13.400 12.200 14.800 13.000 ;
        RECT 13.400 10.600 14.000 13.000 ;
        RECT 11.600 10.600 14.000 11.200 ;
        RECT 11.600 6.800 12.200 11.200 ;
        RECT 11.000 6.600 11.800 7.400 ;
        RECT 1.200 6.800 12.200 7.400 ;
        RECT 5.400 3.800 6.000 7.400 ;
        RECT 5.200 3.800 6.000 4.600 ;
        RECT 4.200 6.800 5.000 7.600 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        RECT 2.600 8.400 3.400 9.200 ;
        RECT 6.800 8.600 7.600 9.400 ;
        RECT 2.600 8.600 7.600 9.200 ;
    END
  END D
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 2.000 -0.600 2.800 5.200 ;
        RECT -0.400 -0.600 19.600 0.600 ;
        RECT 16.400 -0.600 17.200 5.000 ;
        RECT 10.800 -0.600 11.600 3.200 ;
        RECT 7.400 -0.600 8.400 3.200 ;
    END
  END gnd
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 2.000 11.000 2.800 20.600 ;
        RECT -0.400 19.400 19.600 20.600 ;
        RECT 16.400 10.800 17.200 20.600 ;
        RECT 10.800 14.800 11.600 20.600 ;
        RECT 7.600 14.800 8.400 20.600 ;
    END
  END vdd
  OBS 
      LAYER metal2 ;
        RECT 0.400 5.200 1.200 10.800 ;
        RECT 3.600 3.200 4.400 14.800 ;
        RECT 13.200 3.200 14.000 14.800 ;
      LAYER metal1 ;
        RECT 0.400 1.200 1.200 6.000 ;
        RECT 3.600 14.000 4.400 15.400 ;
        RECT 3.600 14.800 5.600 15.400 ;
        RECT 4.800 14.800 5.600 18.800 ;
        RECT 4.800 1.200 5.600 3.200 ;
        RECT 3.600 2.600 5.600 3.200 ;
        RECT 3.600 2.600 4.400 4.000 ;
        RECT 3.600 11.400 9.000 12.000 ;
        RECT 3.600 11.400 4.400 12.200 ;
        RECT 8.200 11.400 9.000 12.200 ;
        RECT 9.200 1.200 10.000 3.200 ;
        RECT 9.200 1.200 9.800 4.400 ;
        RECT 7.000 3.800 9.800 4.400 ;
        RECT 7.000 3.800 7.800 4.600 ;
        RECT 7.000 13.400 7.800 14.200 ;
        RECT 9.800 13.400 10.600 14.200 ;
        RECT 7.000 13.600 10.600 14.200 ;
        RECT 9.200 13.600 9.800 18.800 ;
        RECT 9.200 14.800 10.000 18.800 ;
        RECT 0.400 10.000 6.200 10.400 ;
        RECT 0.400 9.800 6.000 10.400 ;
        RECT 5.400 10.200 10.200 10.800 ;
        RECT 9.600 10.200 10.200 12.600 ;
        RECT 11.000 11.800 11.800 12.600 ;
        RECT 9.600 12.000 11.800 12.600 ;
        RECT 0.400 9.800 1.200 18.800 ;
        RECT 13.200 14.000 14.000 14.800 ;
        RECT 13.400 14.800 14.600 18.800 ;
        RECT 13.400 1.200 14.600 3.200 ;
        RECT 13.200 2.600 14.000 4.000 ;
        RECT 13.200 8.000 14.000 8.800 ;
        RECT 13.200 8.200 17.000 8.800 ;
        RECT 16.200 8.200 17.000 9.000 ;
      LAYER via1 ;
        RECT 0.600 10.200 1.000 10.600 ;
        RECT 0.600 5.400 1.000 5.800 ;
        RECT 3.800 14.200 4.200 14.600 ;
        RECT 3.800 11.600 4.200 12.000 ;
        RECT 3.800 3.400 4.200 3.800 ;
        RECT 13.400 14.200 13.800 14.600 ;
        RECT 13.400 8.200 13.800 8.600 ;
        RECT 13.400 3.400 13.800 3.800 ;
  END 
END DFFPOSX1

MACRO FAX1
  CLASS  CORE ;
  FOREIGN FAX1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 24.000 BY 20.000 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN YC
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        RECT 22.800 1.200 23.600 3.200 ;
        RECT 22.800 14.800 23.600 18.800 ;
        RECT 23.000 1.200 23.600 18.800 ;
        RECT 22.800 6.600 23.600 7.400 ;
    END
  END YC
  PIN YS
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        RECT 19.600 1.200 20.400 3.200 ;
        RECT 20.800 4.600 22.000 5.400 ;
        RECT 19.400 9.200 21.400 9.800 ;
        RECT 20.800 3.800 21.400 9.800 ;
        RECT 19.800 3.800 21.400 4.400 ;
        RECT 19.600 14.800 20.400 18.800 ;
        RECT 19.800 1.200 20.400 4.400 ;
        RECT 19.400 9.200 20.000 15.400 ;
    END
  END YS
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        RECT 0.600 6.000 2.000 6.600 ;
        RECT 17.800 6.800 18.600 7.600 ;
        RECT 17.800 5.600 18.400 7.600 ;
        RECT 7.400 5.600 18.400 6.200 ;
        RECT 0.600 6.000 8.200 6.400 ;
        RECT 1.200 5.800 18.400 6.200 ;
        RECT 0.400 6.600 1.200 7.400 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        RECT 2.200 7.200 2.800 9.400 ;
        RECT 16.000 6.800 16.800 7.600 ;
        RECT 9.400 6.800 16.800 7.400 ;
        RECT 2.200 7.200 10.200 7.600 ;
        RECT 2.800 7.000 16.800 7.400 ;
        RECT 5.800 7.000 6.600 7.800 ;
        RECT 2.200 7.200 3.600 7.800 ;
        RECT 2.000 8.600 2.800 9.400 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        RECT 3.600 8.600 5.200 9.400 ;
        RECT 14.400 8.000 15.200 8.800 ;
        RECT 10.400 8.200 15.200 8.800 ;
        RECT 3.600 8.600 11.800 9.000 ;
        RECT 3.600 8.600 11.000 9.200 ;
    END
  END C
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 2.000 -0.600 2.800 4.000 ;
        RECT -0.400 -0.600 24.400 0.600 ;
        RECT 21.200 -0.600 22.000 3.200 ;
        RECT 18.000 -0.600 18.800 5.000 ;
        RECT 11.000 -0.600 11.800 3.800 ;
        RECT 7.800 -0.600 8.600 4.800 ;
    END
  END gnd
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 2.000 12.000 2.800 20.600 ;
        RECT -0.400 19.400 24.400 20.600 ;
        RECT 21.200 14.800 22.000 20.600 ;
        RECT 18.000 9.200 18.800 20.600 ;
        RECT 11.000 12.800 11.800 20.600 ;
        RECT 7.800 10.800 8.600 20.600 ;
    END
  END vdd
  OBS 
      LAYER metal2 ;
        RECT 14.400 4.200 15.200 5.000 ;
        RECT 14.600 7.800 20.200 8.400 ;
        RECT 19.400 7.800 20.200 8.600 ;
        RECT 14.600 4.200 15.200 10.200 ;
        RECT 14.400 9.400 15.200 10.200 ;
        RECT 5.200 4.400 6.000 5.200 ;
        RECT 12.000 9.600 12.800 11.400 ;
        RECT 20.800 10.600 21.600 11.400 ;
        RECT 5.200 10.800 21.600 11.400 ;
        RECT 5.400 4.400 6.000 11.600 ;
        RECT 5.200 10.800 6.000 11.600 ;
      LAYER metal1 ;
        RECT 0.400 10.800 4.400 11.400 ;
        RECT 0.400 10.800 1.200 18.800 ;
        RECT 3.600 10.800 4.400 18.800 ;
        RECT 0.400 1.200 1.200 5.200 ;
        RECT 3.600 1.200 4.400 5.200 ;
        RECT 0.400 4.600 4.400 5.200 ;
        RECT 5.200 10.800 6.000 18.800 ;
        RECT 5.200 1.200 6.000 5.200 ;
        RECT 9.400 11.600 13.400 12.200 ;
        RECT 9.400 10.800 10.200 18.800 ;
        RECT 12.600 11.600 13.400 18.800 ;
        RECT 9.400 1.200 10.200 5.000 ;
        RECT 12.600 1.200 13.400 5.000 ;
        RECT 9.400 4.400 13.400 5.000 ;
        RECT 12.800 9.400 13.600 10.200 ;
        RECT 12.000 9.600 12.800 10.400 ;
        RECT 14.400 9.400 15.200 18.800 ;
        RECT 14.200 10.200 15.200 18.800 ;
        RECT 14.200 1.200 15.200 4.200 ;
        RECT 14.400 1.200 15.200 5.000 ;
        RECT 19.400 7.000 20.200 8.600 ;
        RECT 20.800 10.600 22.400 11.400 ;
      LAYER via1 ;
        RECT 5.400 11.000 5.800 11.400 ;
        RECT 5.400 4.600 5.800 5.000 ;
        RECT 12.200 9.800 12.600 10.200 ;
        RECT 14.600 9.600 15.000 10.000 ;
        RECT 14.600 4.400 15.000 4.800 ;
        RECT 19.600 8.000 20.000 8.400 ;
        RECT 21.000 10.800 21.400 11.200 ;
  END 
END FAX1

MACRO HAX1
  CLASS  CORE ;
  FOREIGN HAX1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 16.000 BY 20.000 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN YC
    DIRECTION OUTPUT ;
    PORT
      LAYER metal2 ;
        RECT 4.600 3.200 6.000 4.000 ;
        RECT 5.200 8.400 6.000 9.200 ;
        RECT 5.400 3.200 6.000 9.200 ;
      LAYER via1 ;
        RECT 4.800 3.400 5.200 3.800 ;
        RECT 5.400 8.600 5.800 9.000 ;
      LAYER metal1 ;
        RECT 4.600 1.200 5.400 4.000 ;
        RECT 5.200 8.400 6.000 18.800 ;
    END
  END YC
  PIN YS
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        RECT 13.200 10.600 14.000 11.400 ;
        RECT 14.200 14.800 15.000 18.800 ;
        RECT 14.400 13.600 15.000 18.800 ;
        RECT 13.400 4.000 15.000 4.600 ;
        RECT 14.400 1.200 15.000 4.600 ;
        RECT 13.400 13.600 15.000 14.200 ;
        RECT 14.200 1.200 15.000 3.200 ;
        RECT 13.400 4.000 14.000 14.200 ;
    END
  END YS
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        RECT 0.400 6.000 1.200 7.400 ;
        RECT 10.000 6.600 10.800 7.400 ;
        RECT 8.400 6.600 10.800 7.200 ;
        RECT 0.400 6.000 9.000 6.600 ;
        RECT 0.800 5.800 1.600 6.600 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        RECT 2.200 8.000 3.000 8.600 ;
        RECT 8.400 7.800 9.200 8.600 ;
        RECT 7.200 7.800 9.200 8.400 ;
        RECT 2.400 7.200 7.800 7.800 ;
        RECT 2.400 7.200 3.200 8.000 ;
        RECT 2.000 8.600 2.800 9.400 ;
    END
  END B
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.400 -0.600 1.200 5.200 ;
        RECT -0.400 -0.600 16.400 0.600 ;
        RECT 12.600 -0.600 13.400 3.200 ;
        RECT 6.200 -0.600 7.000 5.000 ;
    END
  END gnd
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 2.000 15.200 2.800 20.600 ;
        RECT -0.400 19.400 16.400 20.600 ;
        RECT 12.600 14.800 13.400 20.600 ;
        RECT 11.000 10.800 11.800 20.600 ;
        RECT 6.800 14.800 7.600 20.600 ;
    END
  END vdd
  OBS 
      LAYER metal2 ;
        RECT 3.800 4.600 4.600 5.400 ;
        RECT 3.800 4.600 4.400 9.200 ;
        RECT 3.800 8.400 4.600 9.200 ;
      LAYER metal1 ;
        RECT 3.800 8.400 4.600 9.200 ;
        RECT 0.600 14.000 4.400 14.600 ;
        RECT 0.600 14.000 1.200 18.800 ;
        RECT 0.400 14.800 1.200 18.800 ;
        RECT 3.800 8.400 4.400 18.800 ;
        RECT 3.600 14.000 4.400 18.800 ;
        RECT 3.000 1.200 3.800 5.200 ;
        RECT 3.800 4.600 5.600 5.400 ;
        RECT 7.800 1.200 11.800 1.800 ;
        RECT 11.000 1.200 11.800 4.800 ;
        RECT 7.800 1.200 8.600 5.200 ;
        RECT 9.400 2.400 10.200 5.200 ;
        RECT 9.600 2.400 10.200 6.000 ;
        RECT 9.600 5.400 12.600 6.000 ;
        RECT 11.400 5.400 12.600 6.200 ;
        RECT 11.400 5.400 12.000 10.200 ;
        RECT 8.600 9.600 12.000 10.200 ;
        RECT 8.600 9.600 9.200 18.800 ;
        RECT 8.400 10.800 9.200 18.800 ;
      LAYER via1 ;
        RECT 4.000 8.600 4.400 9.000 ;
        RECT 4.000 4.800 4.400 5.200 ;
  END 
END HAX1

MACRO INVX1
  CLASS  CORE ;
  FOREIGN INVX1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.200 BY 20.000 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        RECT 0.400 3.800 1.200 5.400 ;
    END
  END A
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.400 -0.600 1.200 3.200 ;
        RECT -0.400 -0.600 3.600 0.600 ;
    END
  END gnd
  PIN Y
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        RECT 2.000 1.200 2.800 18.800 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.400 14.800 1.200 20.600 ;
        RECT -0.400 19.400 3.600 20.600 ;
    END
  END vdd
END INVX1

MACRO INVX2
  CLASS  CORE ;
  FOREIGN INVX2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.200 BY 20.000 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        RECT 0.400 5.800 1.200 7.400 ;
    END
  END A
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.400 -0.600 1.200 5.200 ;
        RECT -0.400 -0.600 3.600 0.600 ;
    END
  END gnd
  PIN Y
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        RECT 2.000 1.200 2.800 18.800 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.400 10.800 1.200 20.600 ;
        RECT -0.400 19.400 3.600 20.600 ;
    END
  END vdd
END INVX2

MACRO INVX4
  CLASS  CORE ;
  FOREIGN INVX4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.800 BY 20.000 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        RECT 0.400 5.800 1.200 7.400 ;
    END
  END A
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.400 -0.600 1.200 5.200 ;
        RECT -0.400 -0.600 5.200 0.600 ;
        RECT 3.600 -0.600 4.400 5.200 ;
    END
  END gnd
  PIN Y
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        RECT 2.000 1.200 2.800 18.800 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.400 10.800 1.200 20.600 ;
        RECT -0.400 19.400 5.200 20.600 ;
        RECT 3.600 10.800 4.400 20.600 ;
    END
  END vdd
END INVX4

MACRO INVX8
  CLASS  CORE ;
  FOREIGN INVX8 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.000 BY 20.000 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        RECT 0.400 5.800 1.200 7.400 ;
    END
  END A
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.400 -0.600 1.200 5.200 ;
        RECT -0.400 -0.600 8.400 0.600 ;
        RECT 6.800 -0.600 7.600 5.200 ;
        RECT 3.600 -0.600 4.400 5.200 ;
    END
  END gnd
  PIN Y
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        RECT 2.000 1.200 2.800 6.600 ;
        RECT 5.200 1.200 6.000 18.800 ;
        RECT 2.000 9.400 6.000 10.200 ;
        RECT 2.000 5.800 6.000 6.600 ;
        RECT 2.000 9.400 2.800 18.800 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.400 10.800 1.200 20.600 ;
        RECT -0.400 19.400 8.400 20.600 ;
        RECT 6.800 10.800 7.600 20.600 ;
        RECT 3.600 10.800 4.400 20.600 ;
    END
  END vdd
END INVX8

MACRO NAND2X1
  CLASS  CORE ;
  FOREIGN NAND2X1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.800 BY 20.000 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        RECT 0.400 5.800 1.200 7.400 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        RECT 3.600 10.600 4.400 12.200 ;
    END
  END B
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.400 -0.600 1.200 5.200 ;
        RECT -0.400 -0.600 5.200 0.600 ;
    END
  END gnd
  PIN Y
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        RECT 2.000 4.600 2.800 18.800 ;
        RECT 2.000 4.600 3.800 5.200 ;
        RECT 3.000 1.200 3.800 5.200 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.400 14.800 1.200 20.600 ;
        RECT -0.400 19.400 5.200 20.600 ;
        RECT 3.600 14.800 4.400 20.600 ;
    END
  END vdd
END NAND2X1

MACRO NAND3X1
  CLASS  CORE ;
  FOREIGN NAND3X1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.400 BY 20.000 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        RECT 0.400 9.800 1.200 11.400 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        RECT 2.000 8.600 3.600 9.400 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        RECT 3.600 11.800 4.400 13.400 ;
    END
  END C
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.400 -0.600 1.200 7.200 ;
        RECT -0.400 -0.600 6.800 0.600 ;
    END
  END gnd
  PIN Y
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        RECT 2.200 14.000 2.800 18.800 ;
        RECT 5.200 14.800 6.000 18.800 ;
        RECT 5.200 10.600 6.000 11.400 ;
        RECT 5.200 6.800 5.800 18.800 ;
        RECT 2.200 14.000 5.800 14.600 ;
        RECT 4.200 6.800 5.800 7.400 ;
        RECT 4.000 1.200 4.800 7.200 ;
        RECT 2.000 14.800 2.800 18.800 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.400 14.800 1.200 20.600 ;
        RECT -0.400 19.400 6.800 20.600 ;
        RECT 3.600 15.200 4.400 20.600 ;
    END
  END vdd
END NAND3X1

MACRO NOR2X1
  CLASS  CORE ;
  FOREIGN NOR2X1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.800 BY 20.000 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        RECT 0.400 3.800 1.200 5.400 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        RECT 3.600 8.600 4.400 10.200 ;
    END
  END B
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.400 -0.600 1.200 3.200 ;
        RECT -0.400 -0.600 5.200 0.600 ;
        RECT 3.600 -0.600 4.400 3.200 ;
    END
  END gnd
  PIN Y
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        RECT 2.000 1.200 2.800 3.200 ;
        RECT 3.000 10.800 3.800 18.800 ;
        RECT 2.000 10.800 3.800 11.600 ;
        RECT 2.200 1.200 2.800 11.600 ;
        RECT 2.000 6.600 2.800 7.400 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.400 10.800 1.200 20.600 ;
        RECT -0.400 19.400 5.200 20.600 ;
    END
  END vdd
END NOR2X1

MACRO OAI21X1
  CLASS  CORE ;
  FOREIGN OAI21X1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.400 BY 20.000 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        RECT 0.400 6.600 1.200 7.400 ;
        RECT 1.200 6.200 2.000 7.200 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        RECT 2.000 7.800 2.800 9.400 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        RECT 4.600 10.800 5.200 13.400 ;
        RECT 5.200 10.600 6.000 11.400 ;
        RECT 4.400 12.600 5.200 13.400 ;
    END
  END C
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 2.000 -0.600 2.800 4.400 ;
        RECT -0.400 -0.600 6.800 0.600 ;
    END
  END gnd
  PIN Y
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        RECT 3.000 10.800 3.800 18.800 ;
        RECT 3.400 6.600 6.000 7.400 ;
        RECT 5.200 1.200 6.000 5.200 ;
        RECT 5.200 1.200 5.800 7.400 ;
        RECT 3.400 6.600 4.000 11.400 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.400 10.800 1.200 20.600 ;
        RECT -0.400 19.400 6.800 20.600 ;
        RECT 4.600 14.800 5.400 20.600 ;
    END
  END vdd
  OBS 
      LAYER metal1 ;
        RECT 0.400 1.200 1.200 5.200 ;
        RECT 3.600 1.200 4.400 5.200 ;
        RECT 0.600 5.000 4.200 5.600 ;
  END 
END OAI21X1

MACRO OAI22X1
  CLASS  CORE ;
  FOREIGN OAI22X1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.000 BY 20.000 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        RECT 0.400 6.600 1.200 7.400 ;
        RECT 1.200 6.200 2.000 7.200 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        RECT 2.000 7.800 2.800 9.400 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        RECT 6.800 6.600 7.600 8.200 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        RECT 5.200 7.800 6.000 9.400 ;
    END
  END D
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 2.000 -0.600 2.800 4.400 ;
        RECT -0.400 -0.600 8.400 0.600 ;
    END
  END gnd
  PIN Y
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        RECT 3.600 6.600 4.200 18.800 ;
        RECT 3.600 6.600 6.000 7.200 ;
        RECT 5.400 2.400 6.000 7.200 ;
        RECT 5.200 2.400 6.000 5.200 ;
        RECT 3.000 10.800 5.000 18.800 ;
        RECT 3.600 6.600 4.400 7.400 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.400 10.800 1.200 20.600 ;
        RECT -0.400 19.400 8.400 20.600 ;
        RECT 6.800 10.800 7.600 20.600 ;
    END
  END vdd
  OBS 
      LAYER metal1 ;
        RECT 3.600 1.200 7.600 1.800 ;
        RECT 0.400 1.200 1.200 5.200 ;
        RECT 3.600 1.200 4.400 5.200 ;
        RECT 6.800 1.200 7.600 5.200 ;
        RECT 0.600 5.000 4.200 5.600 ;
  END 
END OAI22X1

MACRO OR2X1
  CLASS  CORE ;
  FOREIGN OR2X1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.400 BY 20.000 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        RECT 0.400 3.800 1.200 5.400 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        RECT 2.000 6.600 2.800 7.400 ;
        RECT 2.200 5.800 3.600 6.600 ;
    END
  END B
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.400 -0.600 1.200 3.200 ;
        RECT -0.400 -0.600 6.800 0.600 ;
        RECT 3.600 -0.600 4.400 3.200 ;
    END
  END gnd
  PIN Y
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        RECT 5.200 1.200 6.000 3.200 ;
        RECT 5.400 1.200 6.000 14.800 ;
        RECT 4.600 14.800 5.400 18.800 ;
        RECT 4.800 14.200 6.000 14.800 ;
        RECT 5.200 8.600 6.000 9.400 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 3.000 10.800 3.800 20.600 ;
        RECT -0.400 19.400 6.800 20.600 ;
    END
  END vdd
  OBS 
      LAYER metal1 ;
        RECT 2.000 1.200 2.800 3.200 ;
        RECT 2.200 1.200 2.800 4.800 ;
        RECT 2.200 4.200 4.800 4.800 ;
        RECT 4.200 4.200 4.800 7.800 ;
        RECT 3.800 7.200 4.400 10.200 ;
        RECT 3.800 9.400 4.600 10.200 ;
        RECT 0.400 9.600 4.600 10.200 ;
        RECT 0.400 9.600 1.200 18.800 ;
  END 
END OR2X1

MACRO OR2X2
  CLASS  CORE ;
  FOREIGN OR2X2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.400 BY 20.000 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        RECT 0.400 3.800 1.200 5.400 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        RECT 2.000 6.600 3.000 7.400 ;
        RECT 2.400 7.400 3.200 8.200 ;
    END
  END B
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.400 -0.600 1.200 3.200 ;
        RECT -0.400 -0.600 6.800 0.600 ;
        RECT 3.600 -0.600 4.400 4.800 ;
    END
  END gnd
  PIN Y
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        RECT 5.200 1.200 6.000 5.200 ;
        RECT 5.400 1.200 6.000 11.400 ;
        RECT 4.600 10.800 5.400 18.800 ;
        RECT 5.200 8.600 6.000 9.400 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 3.000 10.800 3.800 20.600 ;
        RECT -0.400 19.400 6.800 20.600 ;
    END
  END vdd
  OBS 
      LAYER metal1 ;
        RECT 2.000 1.200 2.800 3.200 ;
        RECT 2.200 1.200 2.800 6.000 ;
        RECT 2.200 5.400 4.600 6.000 ;
        RECT 3.800 9.000 4.600 9.800 ;
        RECT 4.000 5.400 4.600 9.800 ;
        RECT 0.400 9.600 4.400 10.200 ;
        RECT 0.400 9.600 1.200 18.800 ;
  END 
END OR2X2

MACRO TBUFX1
  CLASS  CORE ;
  FOREIGN TBUFX1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.000 BY 20.000 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        RECT 6.000 6.600 7.600 7.400 ;
    END
  END A
  PIN EN
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        RECT 0.400 12.600 2.000 13.400 ;
    END
  END EN
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.400 -0.600 1.200 3.200 ;
        RECT -0.400 -0.600 8.400 0.600 ;
        RECT 6.400 -0.600 7.200 5.200 ;
    END
  END gnd
  PIN Y
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        RECT 3.800 1.200 4.600 5.200 ;
        RECT 3.800 10.800 4.600 18.800 ;
        RECT 4.000 1.200 4.600 18.800 ;
        RECT 3.600 8.600 4.600 9.400 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.400 14.800 1.200 20.600 ;
        RECT -0.400 19.400 8.400 20.600 ;
        RECT 6.400 10.800 7.200 20.600 ;
    END
  END vdd
  OBS 
      LAYER metal1 ;
        RECT 2.000 1.200 2.800 3.200 ;
        RECT 2.600 6.600 3.400 7.400 ;
        RECT 2.600 2.400 3.200 8.000 ;
        RECT 2.400 7.400 3.000 10.600 ;
        RECT 2.600 10.000 3.200 15.400 ;
        RECT 2.000 14.800 2.800 18.800 ;
  END 
END TBUFX1

MACRO TBUFX2
  CLASS  CORE ;
  FOREIGN TBUFX2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.200 BY 20.000 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        RECT 9.000 6.600 10.800 7.400 ;
    END
  END A
  PIN EN
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        RECT 0.400 5.800 1.000 10.200 ;
        RECT 0.400 5.800 1.400 6.600 ;
        RECT 0.400 8.600 1.200 10.200 ;
    END
  END EN
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.400 -0.600 1.200 5.200 ;
        RECT -0.400 -0.600 11.600 0.600 ;
        RECT 8.400 -0.600 9.200 4.600 ;
    END
  END gnd
  PIN Y
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        RECT 5.200 2.400 5.800 17.600 ;
        RECT 5.200 10.800 6.000 17.600 ;
        RECT 5.200 8.600 6.000 9.400 ;
        RECT 5.200 2.400 6.000 5.200 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.400 10.800 1.200 20.600 ;
        RECT -0.400 19.400 11.600 20.600 ;
        RECT 8.400 12.200 9.200 20.600 ;
    END
  END vdd
  OBS 
      LAYER metal1 ;
        RECT 2.000 1.200 2.800 5.200 ;
        RECT 2.000 8.200 2.800 9.000 ;
        RECT 2.000 1.200 2.600 18.800 ;
        RECT 2.000 10.800 2.800 18.800 ;
        RECT 6.800 10.800 10.800 11.600 ;
        RECT 3.600 10.800 4.400 18.800 ;
        RECT 6.800 10.800 7.600 18.800 ;
        RECT 3.600 18.200 7.600 18.800 ;
        RECT 10.000 10.800 10.800 18.800 ;
        RECT 3.600 1.200 7.600 1.800 ;
        RECT 10.000 1.200 10.800 4.600 ;
        RECT 6.800 1.200 7.600 5.800 ;
        RECT 3.600 1.200 4.400 5.200 ;
        RECT 10.200 1.200 10.800 5.800 ;
        RECT 6.800 5.200 10.800 5.800 ;
  END 
END TBUFX2

MACRO XOR2X1
  CLASS  CORE ;
  FOREIGN XOR2X1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.200 BY 20.000 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        RECT 0.400 6.600 2.000 7.400 ;
        RECT 4.000 7.000 4.800 7.800 ;
        RECT 2.000 7.000 4.800 7.600 ;
        RECT 0.400 6.800 2.600 7.400 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        RECT 9.200 6.600 10.800 7.400 ;
    END
  END B
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 2.200 -0.600 3.000 4.600 ;
        RECT -0.400 -0.600 11.600 0.600 ;
        RECT 8.200 -0.600 9.200 4.600 ;
        RECT 2.000 1.200 3.000 4.600 ;
    END
  END gnd
  PIN Y
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        RECT 5.200 8.600 6.000 9.400 ;
        RECT 4.800 10.800 6.400 18.800 ;
        RECT 5.800 1.200 6.400 7.400 ;
        RECT 5.400 6.800 6.000 18.800 ;
        RECT 4.800 1.200 6.400 4.800 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 2.000 12.200 3.000 18.800 ;
        RECT -0.400 19.400 11.600 20.600 ;
        RECT 8.200 12.200 9.200 20.600 ;
        RECT 2.200 12.200 3.000 20.600 ;
    END
  END vdd
  OBS 
      LAYER metal2 ;
        RECT 2.200 5.200 3.000 6.000 ;
        RECT 2.200 5.400 7.800 6.000 ;
        RECT 3.600 5.400 4.400 6.200 ;
        RECT 7.000 5.400 7.800 6.200 ;
        RECT 2.200 5.200 2.800 11.600 ;
        RECT 2.200 10.800 3.000 11.600 ;
        RECT 8.400 5.200 9.200 6.000 ;
        RECT 3.600 6.800 9.200 7.400 ;
        RECT 3.600 6.800 4.200 9.600 ;
        RECT 3.400 8.800 4.200 9.600 ;
        RECT 8.600 5.200 9.200 11.600 ;
        RECT 8.400 10.800 9.200 11.600 ;
      LAYER metal1 ;
        RECT 0.400 10.800 3.000 11.400 ;
        RECT 2.200 10.800 3.000 11.600 ;
        RECT 0.400 10.800 1.200 18.800 ;
        RECT 0.400 1.200 1.200 5.800 ;
        RECT 0.400 5.200 3.000 5.800 ;
        RECT 2.200 5.200 3.000 6.000 ;
        RECT 2.600 8.600 3.400 9.400 ;
        RECT 3.400 8.800 4.200 9.600 ;
        RECT 3.600 5.400 5.200 6.200 ;
        RECT 7.000 5.400 7.800 6.200 ;
        RECT 7.200 5.400 7.800 7.400 ;
        RECT 7.200 6.600 8.000 7.400 ;
        RECT 8.400 10.800 10.800 11.400 ;
        RECT 8.400 10.800 9.200 11.600 ;
        RECT 10.000 10.800 10.800 18.800 ;
        RECT 10.000 1.200 10.800 5.800 ;
        RECT 8.400 5.200 10.800 5.800 ;
        RECT 8.400 5.200 9.200 6.000 ;
      LAYER via1 ;
        RECT 2.400 11.000 2.800 11.400 ;
        RECT 2.400 5.400 2.800 5.800 ;
        RECT 3.600 9.000 4.000 9.400 ;
        RECT 3.800 5.600 4.200 6.000 ;
        RECT 7.200 5.600 7.600 6.000 ;
        RECT 8.600 11.000 9.000 11.400 ;
        RECT 8.600 5.400 9.000 5.800 ;
  END 
END XOR2X1

MACRO MUX2X1
  CLASS  CORE ;
  FOREIGN MUX2X1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.600 BY 20.000 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        RECT 6.800 8.600 7.600 10.200 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        RECT 2.000 7.800 2.800 9.400 ;
    END
  END B
  PIN S
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        RECT 0.400 7.800 1.200 9.400 ;
    END
  END S
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 2.000 -0.600 2.800 5.600 ;
        RECT -0.400 -0.600 10.000 0.600 ;
        RECT 7.200 -0.600 8.000 6.000 ;
    END
  END gnd
  PIN Y
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        RECT 4.600 2.000 5.400 5.600 ;
        RECT 5.600 6.600 7.600 7.400 ;
        RECT 4.600 11.200 6.200 11.800 ;
        RECT 5.600 5.000 6.200 11.800 ;
        RECT 5.400 5.000 6.200 6.000 ;
        RECT 4.600 11.200 5.400 18.800 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 2.000 11.200 2.800 20.600 ;
        RECT -0.400 19.400 10.000 20.600 ;
        RECT 7.200 10.800 8.000 20.600 ;
    END
  END vdd
  OBS 
      LAYER metal1 ;
        RECT 0.400 2.000 1.200 4.000 ;
        RECT 0.400 2.000 1.000 6.800 ;
        RECT 0.400 6.200 4.600 6.800 ;
        RECT 3.600 6.200 4.600 8.000 ;
        RECT 3.600 7.200 5.000 8.000 ;
        RECT 3.600 6.200 4.200 10.600 ;
        RECT 0.400 10.000 4.200 10.600 ;
        RECT 0.400 10.000 1.000 18.000 ;
        RECT 0.400 14.000 1.200 18.000 ;
  END 
END MUX2X1

MACRO XNOR2X1
  CLASS  CORE ;
  FOREIGN XNOR2X1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.200 BY 20.000 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER metal2 ;
        RECT 3.600 5.400 4.400 6.200 ;
        RECT 7.000 5.400 7.800 6.200 ;
        RECT 3.600 5.400 7.800 6.000 ;
      LAYER via1 ;
        RECT 3.800 5.600 4.200 6.000 ;
        RECT 7.200 5.600 7.600 6.000 ;
      LAYER metal1 ;
        RECT 0.400 6.600 2.000 7.400 ;
        RECT 7.200 6.600 8.000 7.400 ;
        RECT 7.200 5.400 7.800 7.400 ;
        RECT 7.000 5.400 7.800 6.200 ;
        RECT 3.600 5.400 5.200 6.200 ;
        RECT 0.400 6.600 3.800 7.200 ;
        RECT 3.200 5.600 3.800 7.200 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        RECT 9.200 6.600 10.800 7.400 ;
    END
  END B
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 2.200 -0.600 3.000 4.600 ;
        RECT -0.400 -0.600 11.600 0.600 ;
        RECT 8.200 -0.600 9.200 4.600 ;
        RECT 2.000 1.200 3.000 4.600 ;
    END
  END gnd
  PIN Y
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        RECT 4.800 1.200 6.400 4.800 ;
        RECT 6.200 8.600 7.600 9.400 ;
        RECT 6.200 8.200 6.800 11.400 ;
        RECT 4.800 10.800 6.400 18.800 ;
        RECT 5.800 1.200 6.400 8.800 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 2.000 12.200 3.000 18.800 ;
        RECT -0.400 19.400 11.600 20.600 ;
        RECT 8.200 12.200 9.200 20.600 ;
        RECT 2.200 12.200 3.000 20.600 ;
    END
  END vdd
  OBS 
      LAYER metal2 ;
        RECT 1.800 5.200 2.600 6.000 ;
        RECT 1.800 5.200 2.400 11.600 ;
        RECT 1.800 10.800 2.600 11.600 ;
        RECT 8.400 5.200 9.200 6.000 ;
        RECT 4.400 6.800 9.200 7.400 ;
        RECT 4.400 6.800 5.200 7.600 ;
        RECT 8.600 5.200 9.200 11.600 ;
        RECT 8.400 10.800 9.200 11.600 ;
      LAYER metal1 ;
        RECT 0.400 1.200 1.200 5.800 ;
        RECT 0.400 5.200 2.600 5.800 ;
        RECT 1.800 5.200 2.600 6.000 ;
        RECT 4.400 6.800 5.200 7.600 ;
        RECT 4.400 6.800 5.000 8.800 ;
        RECT 2.400 8.200 5.000 8.800 ;
        RECT 2.400 8.200 3.200 9.000 ;
        RECT 4.600 9.400 5.400 10.200 ;
        RECT 2.000 9.600 5.400 10.200 ;
        RECT 0.400 10.800 2.600 11.400 ;
        RECT 2.000 9.600 2.600 11.600 ;
        RECT 1.800 10.800 2.600 11.600 ;
        RECT 0.400 10.800 1.200 18.800 ;
        RECT 8.400 10.800 10.800 11.400 ;
        RECT 8.400 10.800 9.200 11.600 ;
        RECT 10.000 10.800 10.800 18.800 ;
        RECT 10.000 1.200 10.800 5.800 ;
        RECT 8.400 5.200 10.800 5.800 ;
        RECT 8.400 5.200 9.200 6.000 ;
      LAYER via1 ;
        RECT 2.000 11.000 2.400 11.400 ;
        RECT 2.000 5.400 2.400 5.800 ;
        RECT 4.600 7.000 5.000 7.400 ;
        RECT 8.600 11.000 9.000 11.400 ;
        RECT 8.600 5.400 9.000 5.800 ;
  END 
END XNOR2X1

MACRO LATCH
  CLASS  CORE ;
  FOREIGN LATCH 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.200 BY 20.000 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        RECT 7.400 7.600 10.800 8.400 ;
        RECT 10.000 1.200 10.800 18.800 ;
    END
  END Q
  PIN CLK
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        RECT 1.200 6.600 2.800 7.400 ;
        RECT 5.800 6.600 6.600 8.200 ;
        RECT 1.200 6.600 6.600 7.200 ;
        RECT 4.400 4.600 5.200 7.200 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        RECT 2.600 9.400 4.400 10.200 ;
        RECT 3.600 9.400 4.400 11.400 ;
    END
  END D
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 2.000 -0.600 2.800 5.200 ;
        RECT -0.400 -0.600 11.600 0.600 ;
        RECT 8.400 -0.600 9.200 5.200 ;
    END
  END gnd
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 2.000 10.800 2.800 20.600 ;
        RECT -0.400 19.400 11.600 20.600 ;
        RECT 8.400 10.800 9.200 20.600 ;
    END
  END vdd
  OBS 
      LAYER metal2 ;
        RECT 0.400 5.200 1.200 10.800 ;
        RECT 5.200 3.200 6.000 14.800 ;
      LAYER metal1 ;
        RECT 0.400 9.800 1.200 18.800 ;
        RECT 0.400 1.200 1.200 6.000 ;
        RECT 0.400 8.000 5.000 8.600 ;
        RECT 0.400 8.000 1.200 8.800 ;
        RECT 4.200 8.000 5.000 8.800 ;
        RECT 5.200 14.000 6.000 18.800 ;
        RECT 5.000 14.800 6.200 18.800 ;
        RECT 5.000 1.200 6.200 3.200 ;
        RECT 5.200 1.200 6.000 4.000 ;
        RECT 5.200 9.400 9.400 10.200 ;
      LAYER via1 ;
        RECT 0.600 10.200 1.000 10.600 ;
        RECT 0.600 8.200 1.000 8.600 ;
        RECT 0.600 5.400 1.000 5.800 ;
        RECT 5.400 14.200 5.800 14.600 ;
        RECT 5.400 9.600 5.800 10.000 ;
        RECT 5.400 3.400 5.800 3.800 ;
  END 
END LATCH

MACRO DFFSR
  CLASS  CORE ;
  FOREIGN DFFSR 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 35.200 BY 20.000 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN Q
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        RECT 32.400 1.200 33.200 5.800 ;
        RECT 32.600 5.000 33.400 11.000 ;
        RECT 32.400 10.200 33.200 18.800 ;
    END
  END Q
  PIN CLK
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        RECT 16.400 4.600 18.000 5.400 ;
    END
  END CLK
  PIN R
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        RECT 1.800 8.800 2.600 9.600 ;
        RECT 1.800 9.000 25.200 9.600 ;
        RECT 24.400 8.400 25.200 9.600 ;
        RECT 6.800 8.600 7.600 9.600 ;
    END
  END R
  PIN S
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        RECT 3.600 10.200 4.400 11.400 ;
        RECT 3.600 10.200 30.600 10.800 ;
        RECT 29.800 10.000 30.600 10.800 ;
        RECT 7.000 10.200 7.800 11.000 ;
    END
  END S
  PIN D
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        RECT 13.200 5.800 14.000 7.400 ;
    END
  END D
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 3.600 -0.600 4.400 5.200 ;
        RECT -0.400 -0.600 35.600 0.600 ;
        RECT 34.000 -0.600 34.800 3.200 ;
        RECT 27.600 -0.600 28.400 5.200 ;
        RECT 16.400 -0.600 17.200 3.200 ;
        RECT 13.200 -0.600 14.000 3.200 ;
    END
  END gnd
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.400 14.800 1.200 20.600 ;
        RECT -0.400 19.400 35.600 20.600 ;
        RECT 34.000 14.800 34.800 20.600 ;
        RECT 30.800 14.800 31.600 20.600 ;
        RECT 27.600 14.800 28.400 20.600 ;
        RECT 24.400 14.800 25.200 20.600 ;
        RECT 16.400 14.800 17.200 20.600 ;
        RECT 13.200 14.800 14.000 20.600 ;
        RECT 6.800 14.800 7.600 20.600 ;
        RECT 3.600 14.800 4.400 20.600 ;
    END
  END vdd
  OBS 
      LAYER metal2 ;
        RECT 8.400 3.200 9.200 16.800 ;
        RECT 10.000 3.200 10.800 16.800 ;
        RECT 11.600 3.200 12.400 14.800 ;
        RECT 14.800 3.200 15.600 14.800 ;
        RECT 18.000 3.200 18.800 14.800 ;
        RECT 19.600 3.200 20.400 16.800 ;
        RECT 21.200 3.200 22.000 16.800 ;
        RECT 22.800 3.200 23.600 16.800 ;
      LAYER metal1 ;
        RECT 6.800 1.200 7.600 5.200 ;
        RECT 5.000 4.400 7.600 5.200 ;
        RECT 5.000 4.400 5.800 6.600 ;
        RECT 2.800 5.800 5.800 6.600 ;
        RECT 8.400 16.000 9.200 18.800 ;
        RECT 0.400 7.200 9.200 8.000 ;
        RECT 0.400 1.200 1.200 14.200 ;
        RECT 0.400 13.600 2.400 14.200 ;
        RECT 1.800 13.600 2.400 15.400 ;
        RECT 2.000 14.800 2.800 18.800 ;
        RECT 8.400 1.200 9.200 4.000 ;
        RECT 10.000 16.000 10.800 18.800 ;
        RECT 5.400 11.600 10.800 12.200 ;
        RECT 10.000 11.400 10.800 12.200 ;
        RECT 4.600 12.000 6.000 12.800 ;
        RECT 10.000 1.200 10.800 4.000 ;
        RECT 11.600 14.000 12.400 18.800 ;
        RECT 11.600 1.200 12.400 4.000 ;
        RECT 14.800 14.000 15.600 18.800 ;
        RECT 13.000 12.600 15.600 13.400 ;
        RECT 11.000 4.600 15.600 5.200 ;
        RECT 14.800 4.600 15.600 5.400 ;
        RECT 11.000 4.600 11.800 8.400 ;
        RECT 9.800 7.600 11.800 8.400 ;
        RECT 14.800 1.200 15.600 4.000 ;
        RECT 18.000 12.600 18.800 18.800 ;
        RECT 15.600 7.600 18.800 8.400 ;
        RECT 18.000 1.200 18.800 4.000 ;
        RECT 14.800 6.000 15.600 6.800 ;
        RECT 14.800 6.200 19.200 6.800 ;
        RECT 18.400 6.200 19.200 7.000 ;
        RECT 19.600 16.000 20.400 18.800 ;
        RECT 11.800 11.400 20.400 12.000 ;
        RECT 19.600 11.400 20.400 12.200 ;
        RECT 2.000 12.200 3.600 13.000 ;
        RECT 3.000 12.200 3.600 14.200 ;
        RECT 6.600 12.800 12.400 13.400 ;
        RECT 11.800 11.400 12.400 13.400 ;
        RECT 3.000 13.400 7.200 14.200 ;
        RECT 5.200 13.400 6.000 18.800 ;
        RECT 19.600 1.200 20.400 4.000 ;
        RECT 21.200 16.000 22.000 18.800 ;
        RECT 21.000 4.600 22.000 5.400 ;
        RECT 21.200 4.600 22.000 8.200 ;
        RECT 21.200 1.200 22.000 4.000 ;
        RECT 22.800 16.000 23.600 18.800 ;
        RECT 22.800 1.200 23.600 4.000 ;
        RECT 21.200 13.400 25.400 14.200 ;
        RECT 26.000 12.600 28.600 13.400 ;
        RECT 26.000 12.600 26.800 18.800 ;
        RECT 24.400 1.200 25.200 5.200 ;
        RECT 24.400 4.400 26.800 5.200 ;
        RECT 26.000 4.400 26.800 6.400 ;
        RECT 26.000 5.800 27.800 6.400 ;
        RECT 27.000 5.800 27.800 8.400 ;
        RECT 27.000 7.600 30.800 8.400 ;
        RECT 30.800 1.200 31.600 7.000 ;
        RECT 31.400 6.400 32.000 9.600 ;
        RECT 22.800 11.400 31.800 12.000 ;
        RECT 22.800 11.400 23.600 12.200 ;
        RECT 31.200 9.000 31.800 14.200 ;
        RECT 29.200 13.600 31.800 14.200 ;
        RECT 29.200 13.600 30.000 18.800 ;
      LAYER via1 ;
        RECT 8.600 16.200 9.000 16.600 ;
        RECT 8.600 7.400 9.000 7.800 ;
        RECT 8.600 3.400 9.000 3.800 ;
        RECT 10.200 16.200 10.600 16.600 ;
        RECT 10.200 11.600 10.600 12.000 ;
        RECT 10.200 3.400 10.600 3.800 ;
        RECT 11.800 14.200 12.200 14.600 ;
        RECT 11.800 3.400 12.200 3.800 ;
        RECT 15.000 14.200 15.400 14.600 ;
        RECT 15.000 12.800 15.400 13.200 ;
        RECT 15.000 6.200 15.400 6.600 ;
        RECT 15.000 3.400 15.400 3.800 ;
        RECT 18.200 14.200 18.600 14.600 ;
        RECT 18.200 7.800 18.600 8.200 ;
        RECT 18.200 3.400 18.600 3.800 ;
        RECT 19.800 16.200 20.200 16.600 ;
        RECT 19.800 11.600 20.200 12.000 ;
        RECT 19.800 3.400 20.200 3.800 ;
        RECT 21.400 16.200 21.800 16.600 ;
        RECT 21.400 13.600 21.800 14.000 ;
        RECT 21.400 3.400 21.800 3.800 ;
        RECT 23.000 16.200 23.400 16.600 ;
        RECT 23.000 11.600 23.400 12.000 ;
        RECT 23.000 3.400 23.400 3.800 ;
  END 
END DFFSR

MACRO CLKBUF1
  CLASS  CORE ;
  FOREIGN CLKBUF1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 14.400 BY 20.000 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        RECT 0.400 6.600 1.200 8.000 ;
        RECT 0.400 7.200 2.200 8.000 ;
    END
  END A
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.400 -0.600 1.200 5.200 ;
        RECT -0.400 -0.600 14.800 0.600 ;
        RECT 13.200 -0.600 14.000 5.200 ;
        RECT 10.000 -0.600 10.800 5.200 ;
        RECT 6.800 -0.600 7.600 5.200 ;
        RECT 3.600 -0.600 4.400 5.200 ;
    END
  END gnd
  PIN Y
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        RECT 11.600 1.200 12.400 6.600 ;
        RECT 11.600 9.400 14.000 10.200 ;
        RECT 13.200 5.800 14.000 10.200 ;
        RECT 11.600 5.800 14.000 6.600 ;
        RECT 11.600 9.400 12.400 18.800 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.400 10.800 1.200 20.600 ;
        RECT -0.400 19.400 14.800 20.600 ;
        RECT 13.200 10.800 14.000 20.600 ;
        RECT 10.000 10.800 10.800 20.600 ;
        RECT 6.800 10.800 7.600 20.600 ;
        RECT 3.600 10.800 4.400 20.600 ;
    END
  END vdd
  OBS 
      LAYER metal1 ;
        RECT 2.000 1.200 2.800 6.600 ;
        RECT 2.000 5.800 3.800 6.600 ;
        RECT 3.000 7.200 5.600 8.000 ;
        RECT 3.000 5.800 3.800 10.200 ;
        RECT 2.000 9.400 3.800 10.200 ;
        RECT 2.000 9.400 2.800 18.800 ;
        RECT 5.200 1.200 6.000 6.600 ;
        RECT 5.200 5.800 7.400 6.600 ;
        RECT 6.600 7.200 9.000 8.000 ;
        RECT 6.600 5.800 7.400 10.200 ;
        RECT 5.200 9.400 7.400 10.200 ;
        RECT 5.200 9.400 6.000 18.800 ;
        RECT 8.400 1.200 9.200 6.600 ;
        RECT 8.400 5.800 10.600 6.600 ;
        RECT 9.800 7.200 12.400 8.000 ;
        RECT 9.800 5.800 10.600 10.200 ;
        RECT 8.400 9.400 10.600 10.200 ;
        RECT 8.400 9.400 9.200 18.800 ;
  END 
END CLKBUF1

MACRO CLKBUF2
  CLASS  CORE ;
  FOREIGN CLKBUF2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 20.800 BY 20.000 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        RECT 0.400 6.600 1.200 8.000 ;
        RECT 0.400 7.200 2.200 8.000 ;
    END
  END A
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.400 -0.600 1.200 5.200 ;
        RECT -0.400 -0.600 21.200 0.600 ;
        RECT 19.600 -0.600 20.400 5.200 ;
        RECT 16.400 -0.600 17.200 5.200 ;
        RECT 13.200 -0.600 14.000 5.200 ;
        RECT 10.000 -0.600 10.800 5.200 ;
        RECT 6.800 -0.600 7.600 5.200 ;
        RECT 3.600 -0.600 4.400 5.200 ;
    END
  END gnd
  PIN Y
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        RECT 18.000 1.200 18.800 6.600 ;
        RECT 18.000 9.400 20.400 10.200 ;
        RECT 19.600 5.800 20.400 10.200 ;
        RECT 18.000 5.800 20.400 6.600 ;
        RECT 18.000 9.400 18.800 18.800 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.400 10.800 1.200 20.600 ;
        RECT -0.400 19.400 21.200 20.600 ;
        RECT 19.600 10.800 20.400 20.600 ;
        RECT 16.400 10.800 17.200 20.600 ;
        RECT 13.200 10.800 14.000 20.600 ;
        RECT 10.000 10.800 10.800 20.600 ;
        RECT 6.800 10.800 7.600 20.600 ;
        RECT 3.600 10.800 4.400 20.600 ;
    END
  END vdd
  OBS 
      LAYER metal1 ;
        RECT 2.000 1.200 2.800 6.600 ;
        RECT 2.000 5.800 3.800 6.600 ;
        RECT 3.000 7.200 5.600 8.000 ;
        RECT 3.000 5.800 3.800 10.200 ;
        RECT 2.000 9.400 3.800 10.200 ;
        RECT 2.000 9.400 2.800 18.800 ;
        RECT 5.200 1.200 6.000 6.600 ;
        RECT 5.200 5.800 7.400 6.600 ;
        RECT 6.600 7.200 9.000 8.000 ;
        RECT 6.600 5.800 7.400 10.200 ;
        RECT 5.200 9.400 7.400 10.200 ;
        RECT 5.200 9.400 6.000 18.800 ;
        RECT 8.400 1.200 9.200 6.600 ;
        RECT 8.400 5.800 10.600 6.600 ;
        RECT 9.800 7.200 12.400 8.000 ;
        RECT 9.800 5.800 10.600 10.200 ;
        RECT 8.400 9.400 10.600 10.200 ;
        RECT 8.400 9.400 9.200 18.800 ;
        RECT 11.600 1.200 12.400 6.600 ;
        RECT 11.600 5.800 14.000 6.600 ;
        RECT 13.200 7.200 15.000 8.000 ;
        RECT 13.200 5.800 14.000 10.200 ;
        RECT 11.600 9.400 14.000 10.200 ;
        RECT 11.600 9.400 12.400 18.800 ;
        RECT 14.800 1.200 15.600 6.600 ;
        RECT 14.800 5.800 16.600 6.600 ;
        RECT 15.800 7.200 18.400 8.000 ;
        RECT 15.800 5.800 16.600 10.200 ;
        RECT 14.800 9.400 16.600 10.200 ;
        RECT 14.800 9.400 15.600 18.800 ;
  END 
END CLKBUF2

MACRO CLKBUF3
  CLASS  CORE ;
  FOREIGN CLKBUF3 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 27.200 BY 20.000 ;
  SYMMETRY X Y  ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    PORT
      LAYER metal1 ;
        RECT 0.400 6.600 1.200 8.000 ;
        RECT 0.400 7.200 2.200 8.000 ;
    END
  END A
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.400 -0.600 1.200 5.200 ;
        RECT -0.400 -0.600 27.600 0.600 ;
        RECT 26.000 -0.600 26.800 5.200 ;
        RECT 22.800 -0.600 23.600 5.200 ;
        RECT 19.600 -0.600 20.400 5.200 ;
        RECT 16.400 -0.600 17.200 5.200 ;
        RECT 13.200 -0.600 14.000 5.200 ;
        RECT 10.000 -0.600 10.800 5.200 ;
        RECT 6.800 -0.600 7.600 5.200 ;
        RECT 3.600 -0.600 4.400 5.200 ;
    END
  END gnd
  PIN Y
    DIRECTION OUTPUT ;
    PORT
      LAYER metal1 ;
        RECT 24.400 1.200 25.200 6.600 ;
        RECT 24.400 9.400 26.800 10.200 ;
        RECT 26.000 5.800 26.800 10.200 ;
        RECT 24.400 5.800 26.800 6.600 ;
        RECT 24.400 9.400 25.200 18.800 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.400 10.800 1.200 20.600 ;
        RECT -0.400 19.400 27.600 20.600 ;
        RECT 26.000 10.800 26.800 20.600 ;
        RECT 22.800 10.800 23.600 20.600 ;
        RECT 19.600 10.800 20.400 20.600 ;
        RECT 16.400 10.800 17.200 20.600 ;
        RECT 13.200 10.800 14.000 20.600 ;
        RECT 10.000 10.800 10.800 20.600 ;
        RECT 6.800 10.800 7.600 20.600 ;
        RECT 3.600 10.800 4.400 20.600 ;
    END
  END vdd
  OBS 
      LAYER metal1 ;
        RECT 2.000 1.200 2.800 6.600 ;
        RECT 2.000 5.800 3.800 6.600 ;
        RECT 3.000 7.200 5.600 8.000 ;
        RECT 3.000 5.800 3.800 10.200 ;
        RECT 2.000 9.400 3.800 10.200 ;
        RECT 2.000 9.400 2.800 18.800 ;
        RECT 5.200 1.200 6.000 6.600 ;
        RECT 5.200 5.800 7.400 6.600 ;
        RECT 6.600 7.200 9.000 8.000 ;
        RECT 6.600 5.800 7.400 10.200 ;
        RECT 5.200 9.400 7.400 10.200 ;
        RECT 5.200 9.400 6.000 18.800 ;
        RECT 8.400 1.200 9.200 6.600 ;
        RECT 8.400 5.800 10.600 6.600 ;
        RECT 9.800 7.200 12.400 8.000 ;
        RECT 9.800 5.800 10.600 10.200 ;
        RECT 8.400 9.400 10.600 10.200 ;
        RECT 8.400 9.400 9.200 18.800 ;
        RECT 11.600 1.200 12.400 6.600 ;
        RECT 11.600 5.800 14.000 6.600 ;
        RECT 13.200 7.200 15.000 8.000 ;
        RECT 13.200 5.800 14.000 10.200 ;
        RECT 11.600 9.400 14.000 10.200 ;
        RECT 11.600 9.400 12.400 18.800 ;
        RECT 14.800 1.200 15.600 6.600 ;
        RECT 14.800 5.800 16.600 6.600 ;
        RECT 15.800 7.200 18.400 8.000 ;
        RECT 15.800 5.800 16.600 10.200 ;
        RECT 14.800 9.400 16.600 10.200 ;
        RECT 14.800 9.400 15.600 18.800 ;
        RECT 18.000 1.200 18.800 6.600 ;
        RECT 18.000 5.800 20.200 6.600 ;
        RECT 19.400 7.200 21.800 8.000 ;
        RECT 19.400 5.800 20.200 10.200 ;
        RECT 18.000 9.400 20.200 10.200 ;
        RECT 18.000 9.400 18.800 18.800 ;
        RECT 21.200 1.200 22.000 6.600 ;
        RECT 21.200 5.800 23.400 6.600 ;
        RECT 22.600 7.200 25.200 8.000 ;
        RECT 22.600 5.800 23.400 10.200 ;
        RECT 21.200 9.400 23.400 10.200 ;
        RECT 21.200 9.400 22.000 18.800 ;
  END 
END CLKBUF3

MACRO PADFC
  CLASS  ENDCAP TOPLEFT ;
  FOREIGN PADFC 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 300.000 BY 300.000 ;
  SYMMETRY X Y R90  ;
  SITE corner ;
  OBS 
      LAYER metal4 ;
        RECT 0.600 0.600 299.400 299.400 ;
      LAYER metal3 ;
        RECT 0.600 0.600 299.400 299.400 ;
      LAYER metal2 ;
        RECT 98.000 0.000 170.400 299.400 ;
        RECT 174.800 0.000 195.800 299.400 ;
        RECT 202.200 0.000 223.200 299.400 ;
        RECT 227.600 0.000 300.000 72.400 ;
        RECT 0.600 76.800 300.000 97.800 ;
        RECT 0.600 104.000 300.000 125.200 ;
        RECT 0.600 129.600 300.000 202.000 ;
        RECT 0.600 0.600 299.400 299.400 ;
      LAYER metal1 ;
        RECT 98.000 0.000 195.800 299.400 ;
        RECT 202.200 0.000 300.000 97.800 ;
        RECT 0.600 104.000 300.000 202.000 ;
        RECT 0.600 0.600 299.400 299.400 ;
  END 
END PADFC

MACRO PADGND
  CLASS  PAD ;
  FOREIGN PADGND 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 90.000 BY 300.000 ;
  SYMMETRY R90  ;
  SITE IO ;
  PIN YPAD
    DIRECTION OUTPUT ;
    PORT
      LAYER metal4 ;
        RECT 37.400 254.800 51.200 269.800 ;
    END
  END YPAD
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      CLASS CORE ;
      LAYER metal1 ;
        RECT 34.800 0.000 54.800 0.800 ;
    END
  END gnd
  OBS 
      LAYER metal4 ;
        RECT 0.600 0.600 89.400 253.000 ;
        RECT 0.600 271.600 89.400 299.000 ;
        RECT 0.600 0.600 35.600 299.400 ;
        RECT 53.000 0.600 89.400 299.400 ;
      LAYER metal3 ;
        RECT 0.600 0.600 89.400 299.400 ;
      LAYER metal2 ;
        RECT 0.000 0.000 90.000 72.400 ;
        RECT 0.600 76.600 89.600 97.800 ;
        RECT 0.000 76.800 90.000 97.800 ;
        RECT 0.000 104.200 90.000 125.200 ;
        RECT 0.000 129.600 90.000 202.000 ;
        RECT 0.600 0.000 89.400 299.400 ;
        RECT 6.000 0.000 84.000 300.000 ;
      LAYER metal1 ;
        RECT 0.000 0.000 34.200 97.800 ;
        RECT 55.600 0.000 90.000 97.800 ;
        RECT 0.000 104.200 90.000 202.000 ;
        RECT 0.600 1.800 89.400 299.400 ;
        RECT 6.000 1.800 84.000 300.000 ;
  END 
END PADGND

MACRO PADVDD
  CLASS  PAD ;
  FOREIGN PADVDD 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 90.000 BY 300.000 ;
  SYMMETRY R90  ;
  SITE IO ;
  PIN YPAD
    DIRECTION OUTPUT ;
    PORT
      LAYER metal4 ;
        RECT 42.200 266.000 44.400 268.400 ;
    END
  END YPAD
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      CLASS CORE ;
      LAYER metal1 ;
        RECT 35.400 0.000 54.600 0.800 ;
    END
  END vdd
  OBS 
      LAYER metal4 ;
        RECT 0.600 0.600 89.400 264.200 ;
        RECT 0.600 270.200 89.400 299.000 ;
        RECT 0.600 0.600 40.400 299.400 ;
        RECT 46.200 0.600 89.400 299.400 ;
      LAYER metal3 ;
        RECT 0.600 0.600 89.400 299.400 ;
      LAYER metal2 ;
        RECT 0.000 0.000 34.400 72.400 ;
        RECT 35.400 0.000 54.600 300.000 ;
        RECT 55.600 0.000 90.000 72.400 ;
        RECT 0.000 76.800 90.000 97.800 ;
        RECT 0.000 104.200 90.000 125.200 ;
        RECT 0.000 129.600 90.000 202.000 ;
        RECT 0.600 1.800 89.400 299.400 ;
        RECT 6.000 1.800 84.000 300.000 ;
      LAYER metal1 ;
        RECT 0.000 0.000 34.400 97.800 ;
        RECT 55.600 0.000 90.000 97.800 ;
        RECT 0.000 104.200 90.000 202.000 ;
        RECT 0.600 1.800 89.400 299.400 ;
        RECT 6.000 1.800 84.000 300.000 ;
  END 
END PADVDD

MACRO PADINC
  CLASS  PAD ;
  FOREIGN PADINC 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 90.000 BY 300.000 ;
  SYMMETRY R90  ;
  SITE IO ;
  PIN YPAD
    DIRECTION OUTPUT ;
    PORT
      LAYER metal4 ;
        RECT 42.200 266.000 44.400 268.400 ;
    END
  END YPAD
  PIN DI
    DIRECTION OUTPUT ;
    PORT
      LAYER metal2 ;
        RECT 82.200 -0.400 83.000 0.400 ;
        RECT 81.600 0.000 83.400 0.400 ;
    END
  END DI
  OBS 
      LAYER metal4 ;
        RECT 0.600 0.600 89.400 264.200 ;
        RECT 0.600 270.200 89.400 299.000 ;
        RECT 0.600 0.600 40.400 299.400 ;
        RECT 46.200 0.600 89.400 299.400 ;
      LAYER metal3 ;
        RECT 0.600 0.600 80.600 299.400 ;
        RECT 84.400 0.600 89.400 299.400 ;
        RECT 0.600 1.400 89.400 299.400 ;
      LAYER metal2 ;
        RECT 0.000 0.000 34.400 72.400 ;
        RECT 35.400 0.000 54.600 300.000 ;
        RECT 55.600 0.000 78.200 300.000 ;
        RECT 79.000 0.000 80.800 300.000 ;
        RECT 0.000 0.600 80.800 72.400 ;
        RECT 84.200 0.000 90.000 72.400 ;
        RECT 0.000 76.800 90.000 97.800 ;
        RECT 0.000 104.200 90.000 125.200 ;
        RECT 0.000 129.600 90.000 202.000 ;
        RECT 0.600 1.400 89.400 299.400 ;
        RECT 6.000 1.400 84.000 300.000 ;
      LAYER metal1 ;
        RECT 0.000 0.000 90.000 97.800 ;
        RECT 0.000 104.200 90.000 202.000 ;
        RECT 0.600 0.000 89.400 299.400 ;
        RECT 6.000 0.000 84.000 300.000 ;
  END 
END PADINC

MACRO PADINOUT
  CLASS  PAD ;
  FOREIGN PADINOUT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 90.000 BY 300.000 ;
  SYMMETRY R90  ;
  SITE IO ;
  PIN YPAD
    DIRECTION OUTPUT ;
    PORT
      LAYER metal4 ;
        RECT 42.200 266.000 44.400 268.400 ;
    END
  END YPAD
  PIN DO
    DIRECTION INPUT ;
    PORT
      LAYER metal2 ;
        RECT 8.200 -0.400 9.000 0.400 ;
        RECT 7.600 0.000 9.400 0.400 ;
    END
  END DO
  PIN DI
    DIRECTION OUTPUT ;
    PORT
      LAYER metal2 ;
        RECT 82.200 -0.400 83.000 0.400 ;
        RECT 81.600 0.000 83.400 0.400 ;
    END
  END DI
  PIN OEN
    DIRECTION INPUT ;
    PORT
      LAYER metal2 ;
        RECT 2.600 -0.400 3.400 0.400 ;
        RECT 2.200 0.000 4.000 0.400 ;
    END
  END OEN
  OBS 
      LAYER metal4 ;
        RECT 0.600 0.600 89.400 264.200 ;
        RECT 0.600 270.200 89.400 299.000 ;
        RECT 0.600 0.600 40.400 299.400 ;
        RECT 46.200 0.600 89.400 299.400 ;
      LAYER metal3 ;
        RECT 0.600 0.600 1.200 299.400 ;
        RECT 5.000 0.600 6.600 299.400 ;
        RECT 10.400 0.600 80.600 299.400 ;
        RECT 84.400 0.600 89.400 299.400 ;
        RECT 0.600 1.400 89.400 299.400 ;
      LAYER metal2 ;
        RECT 10.200 0.000 34.400 300.000 ;
        RECT 35.400 0.000 54.600 300.000 ;
        RECT 55.600 0.000 78.200 300.000 ;
        RECT 0.000 0.000 1.400 72.400 ;
        RECT 4.800 0.000 6.800 299.400 ;
        RECT 79.000 0.000 80.800 300.000 ;
        RECT 10.200 0.600 80.800 300.000 ;
        RECT 84.200 0.000 90.000 72.400 ;
        RECT 0.000 76.800 90.000 97.800 ;
        RECT 0.000 104.200 90.000 125.200 ;
        RECT 0.000 129.600 90.000 202.000 ;
        RECT 0.600 1.400 89.400 299.400 ;
        RECT 6.000 1.400 84.000 300.000 ;
      LAYER metal1 ;
        RECT 0.000 0.000 90.000 97.800 ;
        RECT 0.000 104.200 90.000 202.000 ;
        RECT 0.600 0.000 89.400 299.400 ;
        RECT 6.000 0.000 84.000 300.000 ;
  END 
END PADINOUT

MACRO PADNC
  CLASS  PAD ;
  FOREIGN PADNC 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 90.000 BY 300.000 ;
  SYMMETRY R90  ;
  SITE IO ;
  OBS 
      LAYER metal4 ;
        RECT 0.600 0.600 89.400 299.400 ;
      LAYER metal3 ;
        RECT 0.600 0.600 89.400 299.400 ;
      LAYER metal2 ;
        RECT 0.000 0.000 90.000 72.400 ;
        RECT 0.000 76.800 90.000 97.800 ;
        RECT 0.000 104.200 90.000 125.200 ;
        RECT 0.000 129.600 90.000 202.000 ;
        RECT 0.600 0.000 89.400 299.400 ;
      LAYER metal1 ;
        RECT 0.000 0.000 90.000 97.800 ;
        RECT 0.000 104.200 90.000 202.000 ;
        RECT 0.600 0.000 89.400 299.400 ;
  END 
END PADNC

MACRO PADOUT
  CLASS  PAD ;
  FOREIGN PADOUT 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SIZE 90.000 BY 300.000 ;
  SYMMETRY R90  ;
  SITE IO ;
  PIN YPAD
    DIRECTION OUTPUT ;
    PORT
      LAYER metal4 ;
        RECT 42.200 266.000 44.400 268.400 ;
    END
  END YPAD
  PIN DO
    DIRECTION INPUT ;
    PORT
      LAYER metal2 ;
        RECT 8.200 -0.400 9.000 0.400 ;
        RECT 7.600 0.000 9.400 0.400 ;
    END
  END DO
  OBS 
      LAYER metal4 ;
        RECT 0.600 0.600 89.400 264.200 ;
        RECT 0.600 270.200 89.400 299.000 ;
        RECT 0.600 0.600 40.400 299.400 ;
        RECT 46.200 0.600 89.400 299.400 ;
      LAYER metal3 ;
        RECT 0.600 0.600 6.600 299.400 ;
        RECT 10.400 0.600 89.400 299.400 ;
        RECT 0.600 1.400 89.400 299.400 ;
      LAYER metal2 ;
        RECT 0.000 0.000 1.400 72.400 ;
        RECT 2.200 0.000 4.000 299.400 ;
        RECT 4.800 0.000 6.800 299.400 ;
        RECT 10.200 0.000 34.400 300.000 ;
        RECT 35.400 0.000 54.600 300.000 ;
        RECT 55.600 0.000 78.200 300.000 ;
        RECT 79.000 0.000 80.800 300.000 ;
        RECT 81.600 0.000 83.400 300.000 ;
        RECT 0.000 0.600 6.800 72.400 ;
        RECT 10.200 0.600 90.000 72.400 ;
        RECT 84.200 0.000 90.000 72.400 ;
        RECT 0.000 76.800 90.000 97.800 ;
        RECT 0.000 104.200 90.000 125.200 ;
        RECT 0.000 129.600 90.000 202.000 ;
        RECT 0.600 1.400 89.400 299.400 ;
        RECT 6.000 1.400 84.000 300.000 ;
      LAYER metal1 ;
        RECT 0.000 0.000 90.000 97.800 ;
        RECT 0.000 104.200 90.000 202.000 ;
        RECT 0.600 0.000 89.400 299.400 ;
        RECT 6.000 0.000 84.000 300.000 ;
  END 
END PADOUT

END LIBRARY
